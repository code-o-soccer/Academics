`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:32:03 09/08/2019 
// Design Name: 
// Module Name:    barrel 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module barrel(
    input [7:0]inp_,
    input [2:0]shamt,
    input dir,
    output [7:0]out_
    );
	

endmodule
